module synchronizer #(parameter WIDTH = 1) (
                                            input [WIDTH-1:0]  async_signal,
                                            input              clk,
                                            output [WIDTH-1:0] sync_signal
                                            );
endmodule
