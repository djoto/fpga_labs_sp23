module edge_detector #(
                       parameter WIDTH = 1
                       )(
                         input              clk,
                         input [WIDTH-1:0]  signal_in,
                         output [WIDTH-1:0] edge_detect_pulse
                         );
endmodule
